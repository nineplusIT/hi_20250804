`timescale 1ns / 1ps

module tb_SN74_283();

// Port declarations

// DUT

// stimulus

endmodule


