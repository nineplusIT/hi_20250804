`timescale 1ns / 1ps

module tb_traffic_signal_fsm();
  // Port declaration
  
  // internal parameter
  parameter clk_period = 10;

  // DUT
  
  // Reset sequence
  
  // Clock generation
  
  // Stimulus

endmodule
